`include "global.vh"
module DATA_MEMORY
(
    input wire [0:0] SYS_clk,
    input wire [0:0] SYS_reset,

    input wire [1:0]  MEM_write_length,
    input wire [1:0]  MEM_read_length,
    input wire        MEM_read_signed,
    input wire [31:0] MEM_write_data,
    input wire [31:0] MEM_write_address,

    input wire [31:0]  MEM_read_address,

    output reg [31:0] MEM_read_data,
);
    always @(*) 
    begin
        MEM_read_data[31:0]   = {data[MEM_read_address+3],data[MEM_read_address+2], data[MEM_read_address+1], data[MEM_read_address]};
        
        if (MEM_read_length == 2'b01)
        begin
            if (MEM_read_signed)
                MEM_read_data = { {24{data[MEM_read_address][7]}}  , data[MEM_read_address]};
            else 
                MEM_read_data = { {24{1'b0}}  , data[MEM_read_address]};
        end

        else if (MEM_read_length == 2'b10)
        begin
            if (MEM_read_signed)
                MEM_read_data = { {16{data[MEM_read_address + 1][7]}}  , data[MEM_read_address+1], data[MEM_read_address]};
            else 
                MEM_read_data = { {16{1'b0}}  ,                             data[MEM_read_address+1], data[MEM_read_address]};
        end
    end

    integer i;
    always @(posedge SYS_clk) 
    begin
        if (SYS_reset)
        begin
            //TODO Kieungan: initialize the memory in the start of
            $readmemh("C:/Users/tuankiet/Desktop/RISC-v/input_data.txt", data);
        end

        else if (MEM_write_length == 2'b01) //store 1 byte
        begin
            data[MEM_write_address+0] <= MEM_write_data[7:0];
        end

        else if (MEM_write_length == 2'b10) //store half-word
        begin
            data[MEM_write_address+1] <= MEM_write_data[15:8];
            data[MEM_write_address+0] <= MEM_write_data[7:0];
        end

        else if (MEM_write_length == 2'b11) //store word
        begin
            data[MEM_write_address+3] <= MEM_write_data[31:24];
            data[MEM_write_address+2] <= MEM_write_data[23:16];
            data[MEM_write_address+1] <= MEM_write_data[15:8];
            data[MEM_write_address+0] <= MEM_write_data[7:0];
        end
    end

endmodule